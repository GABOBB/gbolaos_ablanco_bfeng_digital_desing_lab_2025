module P1_tb();

endmodule