module P1();

endmodule

